BZh91AY&SY~g1o �_�px��g߰����P�r�ӕ)�$�D����&T�F���z��mM4 &�H=@0F  ��@5=O�M&�j����=A������� s �	������`���`$I�i~��5Oh�1O� ��L�cX 8	*ą`$8�v�$��%�x�ipȒ,4���چ%;����|       "�j�d��d/z:%��SLpRu;)�{�v���W$IX_���=�+IB�s"cE�3A�H���
Ʀ)H�<�`z��w']5ٝ�UUUT*����fffkY���� `�����m��������6�ծt��%��ZMv
�6{&�}�m_���00�.�sAx��\e�s&%#WA*�h@ s��r�������,�fú�e-L"<�.�%s	�Ap�)&�J���)/'�a�A�2�U6ֳ����aBU���36�"�P#a0�рۦ{��ò��*�z)h�CWH��l��x��Ŷ�4 ����T�*RJV�'	��Ɣ���p�L��!!	E+N�I��`��dH�jS!��t5V�,�$�I���"3����]�Z�sz�X�U\:���0�W9z��m�h�Ǫ
j.a��wZ`�k	c�m���~�K[)�p�<�f���T�����j���okۉ�`�Ņy{~mQL������S�����[.C��<u:C  ���I��r� f�Jk4U��Yh���3�Y���$�b�=&�w{-�ٍƢTM���{+ɡ0`�4���/�H�TȁH��&�H1nzdh0P=D�[Ȯ� �ض>U��LV�[�fc[I#X ��"h��|���ʫ1��-���D���Ы�q(�CK '�" ��V���:��gT���_��_Ě5c��H!Hqջ`�ז`��@\�Uðw��e4����E�]ۇ�&A��zLw�	Bd�)�p��4��ގW�l�(k�	�1��%<�n�d�ə�^�h�C�@�2���\D&0踈k�R�-{�"��N�C{�7MÜ�%Ei��yf�����y�FU:m<�����ܑN$��[�